** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/Parametros_Vaf/VTH_tets.sch
**.subckt VTH_tets
N1 Vd Vg GND GND NMOS_ACM w={w} l={l} m=1
V1 Vg GND {Vg}
V2 Vd GND DC({phi_t*0.5})
**** begin user architecture code


* Circuit Parameters
.param vg = 3.0
.param step = 0.01
.param phi_t = 0.0258
.param w = 1.0u
.param l = 1.0u
* Include Models
.model NMOS_ACM nmos_ACM
.model PMOS_ACM pmos_ACM
* OP Parameters & Singals to save
.save all
.save @n1[gm_op]
*Simulations
.dc V1 0 {vg} {step}
.control
pre_osdi NMOS_ACM_2V0.osdi
pre_osdi PMOS_ACM_2V0.osdi
run
let gm_id = deriv(-1*i(V2))/(-1*i(V2))
setplot dc1
gnuplot gm_id
set filetype = ascii
write VTH_sweep.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
