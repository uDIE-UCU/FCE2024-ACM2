** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/Parametros_Vaf/sigma_test.sch
**.subckt sigma_test
N1 Vd Vg GND GND NMOS_ACM w={w} l={l} m=1
E1 Vg GND Vd net1 1000
I0 Vdd Vd {Ibias}
V1 net1 GND {vd}
V2 Vdd GND {vdd}
**** begin user architecture code


* Circuit Parameters
.param vd = 3
.param vdd = 1.2
.param Ibias = 1m
.param step = 0.01
.param w = 5.0u
.param l = 0.18u
* Include Models
.model NMOS_ACM nmos_ACM
.model PMOS_ACM pmos_ACM
* OP Parameters & Singals to save
.save all
.save @n1[gm_op]
.save @n1[gmd_op]
*Simulations
.dc V1 0 {vd} {step}
.control
pre_osdi NMOS_ACM_2V0.osdi
pre_osdi PMOS_ACM_2V0.osdi
run
setplot dc1
plot @n1[gm_op] @n1[gmd_op]
let sigma = @n1[gmd_op]/@n1[gm_op]
set filetype = ascii
write dcsweep.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
