** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/Parametros_Psp/VTH_test_v2.sch
**.subckt VTH_test_v2
V1 Vg GND {Vg}
V2 Vd GND DC({phi_t*0.5})
XM1 Vd Vg GND GND sg13_lv_nmos w={w} l={l} ng=1 m=1
**** begin user architecture code


* Circuit Parameters
.param vg = 3
.param step = 0.01
.param phi_t = 2.4
.param w = 1u
.param l = 100u
* Include Models
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
* OP Parameters & Singals to save
.save all
.save @n.xm1.nsg13_lv_nmos[ide]
.save @n.xm1.nsg13_lv_nmos[gm]
.save @n.xm1.nsg13_lv_nmos[vgs]
.save @n.xm1.nsg13_lv_nmos[vsb]
*Simulations
.dc V1 0 {vg} {step}
.control
run
set filetype = ascii
write dcsweep_v2.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
