** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/Parametros_Psp/n_test.sch
**.subckt n_test
V1 Vs GND {vs}
V2 net1 GND {Vdd}
XM1 Vg Vg Vs GND sg13_lv_nmos w={w} l={l} ng=1 m=1
I0 net1 Vg {is}
**** begin user architecture code


* Circuit Parameters
.param vs = 3
.param step = 0.01
.param Vdd = 1.2
.param is = -0.009377819858216637u
.param w = 1u
.param l = 100u
* Include Models
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
* OP Parameters & Singals to save
.save all
*Simulations
.dc V1 -1 {vs} {step}
.control
run
set filetype = ascii
write dcsweep.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
