** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/Parametros_Psp/VTH_test.sch
**.subckt VTH_test
V1 Vg GND {Vg}
V2 Vd GND DC({phi_t*0.5})
XM1 Vd Vg GND GND sg13_lv_nmos w={w} l={l} ng=1 m=1
**** begin user architecture code


* Circuit Parameters
.param vg = 3
.param step = 0.01
.param phi_t = 0.0258
.param w = 5.0u
.param l = 0.18u
* Include Models
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
* OP Parameters & Singals to save
.save all
*Simulations
.dc V1 0 {vg} {step}
.control
run
setplot dc1
show @n.xm1.nsg13_lv_nmos
let idn = @n.xm1.nsg13_lv_nmos[ids]
let gmn = @n.xm1.nsg13_lv_nmos[gm]
plot ylog abs(idn+i(V2)) idn 0-i(V2)
set filetype = ascii
write dcsweep.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
