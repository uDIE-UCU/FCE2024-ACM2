** sch_path: /workspaces/usm-vlsi-tools/shared_xserver/Parametros_Vaf/zeta_test.sch
**.subckt zeta_test
N1 net1 Vdd GND GND NMOS_ACM w={w} l={l} m=1
V2 Vdd GND {vdd}
Vd Vdd net1 0
.save i(vd)
**** begin user architecture code


* Circuit Parameters
.param vdd = 1.2
.param w = 1.0u
.param l = 1.0u
* Include Models
.model NMOS_ACM nmos_ACM
.model PMOS_ACM pmos_ACM
* OP Parameters & Singals to save
.save all
*Simulations
.op
.control
pre_osdi NMOS_ACM_2V0.osdi
pre_osdi PMOS_ACM_2V0.osdi
run
print i(Vd)
set filetype = ascii
write dcsweep.raw
.endc
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
